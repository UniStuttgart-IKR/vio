--
-- VHDL Package Body riscvio_lib.isa
--
-- Created:
--          by - leylknci.meyer (pc038)
--          at - 19:13:32 04/24/24
--
-- using Mentor Graphics HDL Designer(TM) 2022.3 Built on 14 Jul 2022 at 13:56:12
--
PACKAGE BODY isa IS


    pure function decodeOpc(instruction: std_logic_vector(31 downto 0)) return decode_T is
        variable res: decode_T;
    begin
        res.imm_mode := none;
        case instruction(OPC_RANGE) is
            when OPC_ALU_R => 
                res.imm_mode := none;
                res.me_mode  := holiday;
                res.at_mode  := holiday;
                res.rdst     := to_integer(unsigned(instruction(RD_RANGE)));
                res.rdat     := to_integer(unsigned(instruction(RS1_RANGE)));
                res.rptr     := 0;
                res.raux     := to_integer(unsigned(instruction(RS2_RANGE)));
                case instruction(FUNCT3_RANGE) is
                    when F3_ADD_SUB =>
                        case instruction(FUNCT7_RANGE) is 
                            when F7_ADD_SRL_SLL_XOR_OR_AND_SLT_SLTU =>
                                res.mnemonic := add_r;
                                res.alu_mode := alu_add;
                            when F7_SUB_SRA =>
                                res.mnemonic := sub_r;
                                res.alu_mode := alu_sub;
                            when others =>
                                res.mnemonic := illegal;
                                res.alu_mode := alu_illegal;
                        end case;
                    when (F3_SRL_SRA or F3_MINU_ROR_RORI_ORC_REV) =>
                        res.mnemonic := srl_r when instruction(FUNCT7_RANGE) = F7_ADD_SRL_SLL_XOR_OR_AND_SLT_SLTU else 
                                        sra_i when instruction(FUNCT7_RANGE) = F7_SUB_SRA else 
                                        minu when instruction(FUNCT7_RANGE) = F7_MAX_MAXU_MIN_MINU else 
                                        ror_r when instruction(FUNCT7_RANGE) = F7_CLZ_CTZ_CPOP_SEXT_ROL_ROR else
                                        illegal;
                        res.alu_mode := alu_srl when instruction(FUNCT7_RANGE) = F7_ADD_SRL_SLL_XOR_OR_AND_SLT_SLTU else 
                                        alu_sra when instruction(FUNCT7_RANGE) = F7_SUB_SRA else 
                                        alu_minu when instruction(FUNCT7_RANGE) = F7_MAX_MAXU_MIN_MINU else 
                                        alu_ror when instruction(FUNCT7_RANGE) = F7_CLZ_CTZ_CPOP_SEXT_ROL_ROR else
                                        alu_illegal;
                    when (F3_SLL or F3_ROL_CTZ_CPOP_SEXT) =>
                        res.mnemonic := rol_r when instruction(FUNCT7_RANGE) = F7_CLZ_CTZ_CPOP_SEXT_ROL_ROR else sll_r;
                        res.alu_mode := alu_rol when instruction(FUNCT7_RANGE) = F7_CLZ_CTZ_CPOP_SEXT_ROL_ROR else alu_sll;
                    when F3_SLT =>
                        res.mnemonic := slt_r;
                        res.alu_mode := alu_slt;
                    when F3_SLTU =>
                        res.mnemonic := sltu_r;
                        res.alu_mode := alu_sltu;
                    when (F3_XOR or F3_XNOR_MIN_ZEXT) =>
                        res.mnemonic := xor_r when instruction(FUNCT7_RANGE) = F7_ADD_SRL_SLL_XOR_OR_AND_SLT_SLTU else 
                                        xnor_r when instruction(FUNCT7_RANGE) = F7_ANDN_ORN_XNOR else 
                                        min when instruction(FUNCT7_RANGE) = F7_MAX_MAXU_MIN_MINU else
                                        zext_h when (instruction(FUNCT7_RANGE) = F7_ZEXT and instruction(RS2_RANGE) = F5_CLZ_ZEXT) else 
                                        illegal;
                        res.alu_mode := alu_xor when instruction(FUNCT7_RANGE) = F7_ADD_SRL_SLL_XOR_OR_AND_SLT_SLTU else 
                                        alu_xnor when instruction(FUNCT7_RANGE) = F7_ANDN_ORN_XNOR else 
                                        alu_min when instruction(FUNCT7_RANGE) = F7_MAX_MAXU_MIN_MINU else
                                        alu_zexth when (instruction(FUNCT7_RANGE) = F7_ZEXT and instruction(RS2_RANGE) = F5_CLZ_ZEXT) else 
                                        alu_illegal;
                    when (F3_OR or F3_ORN_MAX) =>
                        res.mnemonic := or_r when instruction(FUNCT7_RANGE) = F7_ADD_SRL_SLL_XOR_OR_AND_SLT_SLTU else 
                                        orn_r when instruction(FUNCT7_RANGE) = F7_ANDN_ORN_XNOR else 
                                        max when instruction(FUNCT7_RANGE) = F7_MAX_MAXU_MIN_MINU else
                                        illegal;
                        res.alu_mode := alu_or when instruction(FUNCT7_RANGE) = F7_ADD_SRL_SLL_XOR_OR_AND_SLT_SLTU else 
                                        alu_orn when instruction(FUNCT7_RANGE) = F7_ANDN_ORN_XNOR else 
                                        alu_max when instruction(FUNCT7_RANGE) = F7_MAX_MAXU_MIN_MINU else
                                        alu_illegal;
                    when F3_AND =>
                        res.mnemonic := and_r when instruction(FUNCT7_RANGE) = F7_ADD_SRL_SLL_XOR_OR_AND_SLT_SLTU else
                                        andn_r when instruction(FUNCT7_RANGE) = F7_ANDN_ORN_XNOR else 
                                        maxu when instruction(FUNCT7_RANGE) = F7_MAX_MAXU_MIN_MINU else
                                        illegal;
                        res.alu_mode := alu_and when instruction(FUNCT7_RANGE) = F7_ADD_SRL_SLL_XOR_OR_AND_SLT_SLTU else
                                        alu_andn when instruction(FUNCT7_RANGE) = F7_ANDN_ORN_XNOR else 
                                        alu_maxu when instruction(FUNCT7_RANGE) = F7_MAX_MAXU_MIN_MINU else
                                        alu_illegal;
                    when others =>
                        res.mnemonic := illegal;
                        res.alu_mode := alu_illegal;
                end case;

            when OPC_ALU_I => 
                res.imm_mode := i_type;
                res.me_mode  := holiday;
                res.at_mode  := holiday;
                res.rdst     := to_integer(unsigned(instruction(RD_RANGE)));
                res.rdat     := to_integer(unsigned(instruction(RS1_RANGE)));
                res.rptr     := 0;
                res.raux     := 0;
                case instruction(FUNCT3_RANGE) is
                    when F3_ADD_SUB =>
                        res.mnemonic := nop when instruction = NOP_INSTR else add_i;
                        res.alu_mode := alu_add;
                    when (F3_SRL_SRA or F3_MINU_ROR_RORI_ORC_REV) =>
                        res.mnemonic := srl_i when instruction(FUNCT7_RANGE) = F7_ADD_SRL_SLL_XOR_OR_AND_SLT_SLTU else
                                        sra_i when instruction(FUNCT7_RANGE) = F7_SUB_SRA else
                                        ror_i when instruction(FUNCT7_RANGE) = F7_CLZ_CTZ_CPOP_SEXT_ROL_ROR else
                                        orcv_b when instruction(FUNCT7_RANGE) = F7_ORC and instruction(RS2_RANGE) = F5_ORC else 
                                        rev8 when instruction(FUNCT7_RANGE) = F7_REV8 and instruction(RS2_RANGE) = F5_REV8 else 
                                        illegal;
                        res.alu_mode := alu_srl when instruction(FUNCT7_RANGE) = F7_ADD_SRL_SLL_XOR_OR_AND_SLT_SLTU else
                                        alu_sra when instruction(FUNCT7_RANGE) = F7_SUB_SRA else
                                        alu_ror when instruction(FUNCT7_RANGE) = F7_CLZ_CTZ_CPOP_SEXT_ROL_ROR else
                                        alu_orcb when instruction(FUNCT7_RANGE) = F7_ORC and instruction(RS2_RANGE) = F5_ORC else 
                                        alu_rev8 when instruction(FUNCT7_RANGE) = F7_REV8 and instruction(RS2_RANGE) = F5_REV8 else 
                                        alu_illegal;
                    when F3_SLT =>
                        res.mnemonic := slt_i;
                        res.alu_mode := alu_slt;
                    when F3_SLTU =>
                        res.mnemonic := sltu_i;
                        res.alu_mode := alu_sltu;
                    when F3_XOR =>
                        res.mnemonic := xor_i;
                        res.alu_mode := alu_xor;
                    when F3_OR =>
                        res.mnemonic := or_i;
                        res.alu_mode := alu_or;
                    when F3_AND =>
                        res.mnemonic := and_i;
                        res.alu_mode := alu_and;
                    when (F3_SLL or F3_ROL_CTZ_CPOP_SEXT) =>
                        if instruction(FUNCT7_RANGE) = F7_ADD_SRL_SLL_XOR_OR_AND_SLT_SLTU then
                            res.mnemonic := sll_i;
                            res.alu_mode := alu_sll;
                        elsif instruction(FUNCT7_RANGE) = F7_CLZ_CTZ_CPOP_SEXT_ROL_ROR then
                            case instruction(RS2_RANGE) is
                                when F5_CLZ_ZEXT => res.mnemonic := clz;
                                                    res.alu_mode := alu_clz;
                                when F5_CTZ =>      res.mnemonic := ctz;
                                                    res.alu_mode := alu_ctz;
                                when F5_CPOP =>     res.mnemonic := cpop;
                                                    res.alu_mode := alu_cpop;
                                when F5_SEXTB =>    res.mnemonic := sext_b;
                                                    res.alu_mode := alu_sextb;
                                when F5_SEXTH =>    res.mnemonic := sext_h;
                                                    res.alu_mode := alu_sexth;
                                when others =>      res.mnemonic := illegal;
                                                    res.alu_mode := alu_illegal;
                            end case;
                        end if;
                    when others =>
                        res.mnemonic := illegal;
                        res.alu_mode := alu_illegal;
                end case;
            when OPC_JAL =>
                res.mnemonic := jal;
                res.alu_mode := alu_illegal;
                res.imm_mode := j_type;
                res.me_mode  := holiday;
                res.at_mode  := holiday;
                res.rdst     := 1 when to_integer(unsigned(instruction(RD_RANGE))) = 1 else 0; --only rix or zero are allowed!
                res.rdat     := 0; 
                res.rptr     := 2; --frame
                res.raux     := 0;
            when OPC_BRANCH =>
                res.alu_mode := alu_add;
                res.imm_mode := b_type;
                res.me_mode  := holiday;
                res.at_mode  := holiday;
                res.rdst     := 0;
                res.rdat     := to_integer(unsigned(instruction(RS1_RANGE)));
                res.rptr     := 0;
                res.raux     := to_integer(unsigned(instruction(RS2_RANGE)));
                case instruction(FUNCT3_RANGE) is
                    when F3_BEQ  => res.mnemonic := beq;
                    when F3_BNE  => res.mnemonic := bne;
                    when F3_BLT  => res.mnemonic := blt;
                    when F3_BGE  => res.mnemonic := bge;
                    when F3_BLTU => res.mnemonic := bltu;
                    when F3_BGEU => res.mnemonic := bgeu;
                    when others =>  res.mnemonic := illegal;
                end case;
            when OPC_LOAD =>
                res.alu_mode := alu_add;
                res.imm_mode := i_type when instruction(FUNCT3_RANGE) /= "111" else none;
                res.me_mode  := load;
                res.at_mode  := holiday;
                res.rdst     := to_integer(unsigned(instruction(RD_RANGE)));
                res.rdat     := to_integer(unsigned(instruction(RS2_RANGE))) when instruction(FUNCT3_RANGE) = "111" else 0;
                res.rptr     := to_integer(unsigned(instruction(RS1_RANGE)));
                res.raux     := 0;
                case instruction(FUNCT3_RANGE) is
                    when F3_BYTE  => res.mnemonic := lb_i;
                    when F3_HALF  => res.mnemonic := lh_i;
                    when F3_WORD  => res.mnemonic := lw_i;
                    when F3_BYTEU => res.mnemonic := lbu_i;
                    when F3_HALFU => res.mnemonic := lhu_i;
                    when F3_REG   => res.mnemonic := illegal;
                    when others =>  res.mnemonic := illegal;
                end case;
            when OPC_STORE =>
                res.alu_mode := alu_add;
                res.imm_mode := s_type when instruction(FUNCT3_RANGE) /= "111" else none;
                res.me_mode  := store;
                res.at_mode  := holiday;
                res.rdst     := 0;
                res.rdat     := to_integer(unsigned(instruction(RD_RANGE))) when instruction(FUNCT3_RANGE) = "111" else 0;
                res.rptr     := to_integer(unsigned(instruction(RS1_RANGE)));
                res.raux     := to_integer(unsigned(instruction(RS2_RANGE)));
                case instruction(FUNCT3_RANGE) is
                    when F3_BYTE  => res.mnemonic := sb_i;
                    when F3_HALF  => res.mnemonic := sh_i;
                    when F3_WORD  => res.mnemonic := sw_i;
                    when F3_REG   => res.mnemonic := illegal;
                    when others =>  res.mnemonic := illegal;
                end case;
            when others =>
                res.mnemonic := illegal;
                res.alu_mode := alu_illegal;
                res.imm_mode := none;
                res.me_mode  := holiday;
                res.at_mode  := holiday;
                res.rdst     := 0;
                res.rdat     := 0;
                res.rptr     := 0;
                res.raux     := 0;
        end case;
        return res;
    end function decodeOpc;

    pure function extractJTypeImm(inst: word_T) return word_T is
        variable res: word_T;
    begin
        res := (0 => '0', others => inst(31));
        res(19 downto 12) := inst(19 downto 12);
        res(11) := inst(20);
        res(10 downto 1) := inst(30 downto 21);
        return res;
    end function extractJTypeImm;


    pure function extractBTypeImm(inst: word_T) return word_T is
        variable res: word_T;
    begin
        res := (0 => '0', others => inst(31));
        res(10 downto 5) := inst(30 downto 25);
        res(11) := inst(7);
        res(4 downto 1) := inst(11 downto 8);
        return res;
    end function extractBTypeImm;

    pure function extractSTypeImm(inst: word_T) return word_T is
        variable res: word_T;
    begin
        res := (others => inst(31));
        res(10 downto 5) := inst(30 downto 25);
        res(4 downto 0) := inst(11 downto 7);
        return res;
    end function extractSTypeImm;

END isa;
