--
-- VHDL Architecture riscvio_lib.ex_reg.behav
--
-- Created:
--          by - surfer.UNKNOWN (SURFER-A0000001)
--          at - 14:00:34 09.05.2024
--
-- using Mentor Graphics HDL Designer(TM) 2021.1 Built on 14 Jan 2021 at 15:11:42
--
ARCHITECTURE behav OF ex_reg IS
BEGIN
      process(clk, res_n) is
    begin
        if res_n = '0' then
        rd_me <= REG_NULL;
        rs1_me <= REG_NULL;
        rs2_me <= REG_NULL;
        ctrl_me <= CTRL_NULL;
        alu_out_me <= (others => '0');
        else
            if clk'event and clk = '1' then
                ctrl_me <= ctrl_ex;

                rs1_me <= rs1_ex;
                rs2_me <= rs2_ex;
                rd_me <= rd_ex;

                alu_out_me <= alu_out_ex_u;
            end if;
        end if;
    end process;

END ARCHITECTURE behav;

