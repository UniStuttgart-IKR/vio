LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY riscvio_lib;
USE riscvio_lib.isa.all;
USE riscvio_lib.pipeline.all;

ENTITY pgu IS
   PORT( 
      imm      : IN     word_T;
      pc       : IN     pc_T;
      pgu_mode : IN     pgu_mode_T;
      raux     : IN     raux_T;
      rdat     : IN     rdat_T;
      rdst_ix  : IN     reg_nbr_T;
      rptr     : IN     rptr_T;
      me_addr  : OUT    mem_addr_T;
      pgu_exc  : OUT    exc_cause_T;
      ptr      : OUT    reg_mem_T
   );

-- Declarations

END pgu ;
