--
-- VHDL Architecture riscvio_lib.alu_mux.behav
--
-- Created:
--          by - leylknci.meyer (pc024)
--          at - 16:42:07 05/22/24
--
-- using Mentor Graphics HDL Designer(TM) 2022.3 Built on 14 Jul 2022 at 13:56:12
--
ARCHITECTURE behav OF alu_a_mux IS
BEGIN
    a <= rdat_dc.val when alu_a_in_sel = DAT else
         rptr_dc.val when alu_a_in_sel = PTRVAL else
         rptr_dc.pi  when alu_a_in_sel = PTRPI else
         rptr_dc.dt  when alu_a_in_sel = PTRDT else
         raux_dc.val;

END ARCHITECTURE behav;

