LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY riscvio_tb IS
-- Declarations

END riscvio_tb ;

