LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY riscvio_soc_tb IS
-- Declarations

END riscvio_soc_tb ;
