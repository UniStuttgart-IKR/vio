LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY riscvio_lib;
USE riscvio_lib.pipeline.all;
USE riscvio_lib.ISA.all;
USE ieee.numeric_std.all;
USE ieee.math_real.all;


ARCHITECTURE struct OF riscvio_soc IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL ac_rack             : boolean;
   SIGNAL ac_raddr            : std_logic_vector(ADDR_WIDTH - 1 DOWNTO 0) := (others => '0');
   SIGNAL ac_rdata            : std_logic_vector(BUS_WIDTH - 1 DOWNTO 0);
   SIGNAL ac_rreq             : boolean                                   := false;
   SIGNAL data_stream_in      : std_logic_vector(7 DOWNTO 0);
   SIGNAL data_stream_in_ack  : std_logic;
   SIGNAL data_stream_in_done : std_logic;
   SIGNAL data_stream_in_stb  : std_logic;
   SIGNAL data_stream_out     : std_logic_vector(7 DOWNTO 0);
   SIGNAL data_stream_out_stb : std_logic;
   SIGNAL dc_rack             : boolean;
   SIGNAL dc_raddr            : std_logic_vector(ADDR_WIDTH - 1 DOWNTO 0) := (others => '0');
   SIGNAL dc_rdata            : std_logic_vector(BUS_WIDTH - 1 DOWNTO 0);
   SIGNAL dc_rreq             : boolean                                   := false;
   SIGNAL dc_wack             : boolean;
   SIGNAL dc_waddr            : std_logic_vector(ADDR_WIDTH - 1 DOWNTO 0) := (others => '0');
   SIGNAL dc_wbyte_ena        : std_logic_vector(BUS_WIDTH/8 - 1 DOWNTO 0);
   SIGNAL dc_wdata            : std_logic_vector(BUS_WIDTH - 1 DOWNTO 0)  := (others => '0');
   SIGNAL dc_wreq             : boolean                                   := false;
   SIGNAL ic_rack             : boolean;
   SIGNAL ic_raddr            : std_logic_vector(ADDR_WIDTH - 1 DOWNTO 0) := (others => '0');
   SIGNAL ic_rdata            : std_logic_vector(BUS_WIDTH - 1 DOWNTO 0);
   SIGNAL ic_rreq             : boolean                                   := false;
   SIGNAL io_dev              : std_logic_vector(11 DOWNTO 0);
   SIGNAL io_ix               : word_T;
   SIGNAL io_mode             : mem_mode_T;
   SIGNAL io_rdata            : word_T;
   SIGNAL io_stall            : std_logic;
   SIGNAL io_wdata            : word_T;


   -- Component Declarations
   COMPONENT int_ram
   PORT (
      ac_raddr     : IN     std_logic_vector (ADDR_WIDTH - 1 DOWNTO 0) := (others => '0');
      ac_rreq      : IN     boolean                                    := false;
      clk          : IN     std_logic;
      dc_raddr     : IN     std_logic_vector (ADDR_WIDTH - 1 DOWNTO 0) := (others => '0');
      dc_rreq      : IN     boolean                                    := false;
      dc_waddr     : IN     std_logic_vector (ADDR_WIDTH - 1 DOWNTO 0) := (others => '0');
      dc_wbyte_ena : IN     std_logic_vector (BUS_WIDTH/8 - 1 DOWNTO 0);
      dc_wdata     : IN     std_logic_vector (BUS_WIDTH - 1 DOWNTO 0)  := (others => '0');
      dc_wreq      : IN     boolean                                    := false;
      ic_raddr     : IN     std_logic_vector (ADDR_WIDTH - 1 DOWNTO 0) := (others => '0');
      ic_rreq      : IN     boolean                                    := false;
      res_n        : IN     std_logic;
      ac_rack      : OUT    boolean;
      ac_rdata     : OUT    std_logic_vector (BUS_WIDTH - 1 DOWNTO 0);
      dc_rack      : OUT    boolean;
      dc_rdata     : OUT    std_logic_vector (BUS_WIDTH - 1 DOWNTO 0);
      dc_wack      : OUT    boolean;
      ic_rack      : OUT    boolean;
      ic_rdata     : OUT    std_logic_vector (BUS_WIDTH - 1 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT io_mux
   PORT (
      clk                 : IN     std_logic ;
      data_stream_in_ack  : IN     std_logic ;
      data_stream_in_done : IN     std_logic ;
      data_stream_out     : IN     std_logic_vector (7 DOWNTO 0);
      data_stream_out_stb : IN     std_logic ;
      io_dev              : IN     std_logic_vector (11 DOWNTO 0);
      io_ix               : IN     word_T ;
      io_mode             : IN     mem_mode_T ;
      io_wdata            : IN     word_T ;
      res_n               : IN     std_logic ;
      data_stream_in      : OUT    std_logic_vector (7 DOWNTO 0);
      data_stream_in_stb  : OUT    std_logic ;
      io_rdata            : OUT    word_T ;
      io_stall            : OUT    std_logic 
   );
   END COMPONENT;
   COMPONENT riscvio
   PORT (
      ac_rack      : IN     boolean ;
      ac_rdata     : IN     buzz_word_T ;
      clk          : IN     std_logic ;
      dc_rack      : IN     boolean ;
      dc_rdata     : IN     buzz_word_T ;
      dc_wack      : IN     boolean ;
      ic_rack      : IN     boolean ;
      ic_rdata     : IN     std_logic_vector (BUS_WIDTH - 1 DOWNTO 0);
      io_rdata     : IN     word_T ;
      io_stall     : IN     std_logic ;
      res_n        : IN     std_logic ;
      ac_raddr     : OUT    std_logic_vector (31 DOWNTO 0);
      ac_rreq      : OUT    boolean ;
      dc_raddr     : OUT    std_logic_vector (31 DOWNTO 0);
      dc_rreq      : OUT    boolean ;
      dc_waddr     : OUT    std_logic_vector (31 DOWNTO 0);
      dc_wbyte_ena : OUT    std_logic_vector (BUS_WIDTH/8 - 1 DOWNTO 0);
      dc_wdata     : OUT    buzz_word_T ;
      dc_wreq      : OUT    boolean ;
      ic_raddr     : OUT    std_logic_vector (ADDR_WIDTH - 1 DOWNTO 0);
      ic_rreq      : OUT    boolean ;
      io_dev       : OUT    std_logic_vector (11 DOWNTO 0);
      io_ix        : OUT    word_T ;
      io_mode      : OUT    mem_mode_T ;
      io_wdata     : OUT    word_T 
   );
   END COMPONENT;
   COMPONENT uart
   GENERIC (
      baud            : positive;
      clock_frequency : positive
   );
   PORT (
      clock               : IN     std_logic;
      data_stream_in      : IN     std_logic_vector (7 DOWNTO 0);
      data_stream_in_stb  : IN     std_logic;
      res_n               : IN     std_logic;
      rx                  : IN     std_logic;
      data_stream_in_ack  : OUT    std_logic;
      data_stream_in_done : OUT    std_logic;
      data_stream_out     : OUT    std_logic_vector (7 DOWNTO 0);
      data_stream_out_stb : OUT    std_logic;
      tx                  : OUT    std_logic
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : int_ram USE ENTITY riscvio_lib.int_ram;
   FOR ALL : io_mux USE ENTITY riscvio_lib.io_mux;
   FOR ALL : riscvio USE ENTITY riscvio_lib.riscvio;
   FOR ALL : uart USE ENTITY riscvio_lib.uart;
   -- pragma synthesis_on


BEGIN

   -- Instance port mappings.
   int_ram_i : int_ram
      PORT MAP (
         clk          => clk,
         res_n        => res_n,
         dc_rreq      => dc_rreq,
         dc_rack      => dc_rack,
         dc_raddr     => dc_raddr,
         dc_rdata     => dc_rdata,
         ac_rreq      => ac_rreq,
         ac_rack      => ac_rack,
         ac_raddr     => ac_raddr,
         ac_rdata     => ac_rdata,
         ic_rreq      => ic_rreq,
         ic_rack      => ic_rack,
         ic_raddr     => ic_raddr,
         ic_rdata     => ic_rdata,
         dc_wreq      => dc_wreq,
         dc_wack      => dc_wack,
         dc_waddr     => dc_waddr,
         dc_wdata     => dc_wdata,
         dc_wbyte_ena => dc_wbyte_ena
      );
   io_mux_i : io_mux
      PORT MAP (
         clk                 => clk,
         data_stream_in_ack  => data_stream_in_ack,
         data_stream_in_done => data_stream_in_done,
         data_stream_out     => data_stream_out,
         data_stream_out_stb => data_stream_out_stb,
         io_dev              => io_dev,
         io_ix               => io_ix,
         io_mode             => io_mode,
         io_wdata            => io_wdata,
         res_n               => res_n,
         data_stream_in      => data_stream_in,
         data_stream_in_stb  => data_stream_in_stb,
         io_rdata            => io_rdata,
         io_stall            => io_stall
      );
   riscvio_i : riscvio
      PORT MAP (
         ac_rack      => ac_rack,
         ac_rdata     => ac_rdata,
         clk          => clk,
         dc_rack      => dc_rack,
         dc_rdata     => dc_rdata,
         dc_wack      => dc_wack,
         ic_rack      => ic_rack,
         ic_rdata     => ic_rdata,
         io_rdata     => io_rdata,
         io_stall     => io_stall,
         res_n        => res_n,
         ac_raddr     => ac_raddr,
         ac_rreq      => ac_rreq,
         dc_raddr     => dc_raddr,
         dc_rreq      => dc_rreq,
         dc_waddr     => dc_waddr,
         dc_wbyte_ena => dc_wbyte_ena,
         dc_wdata     => dc_wdata,
         dc_wreq      => dc_wreq,
         ic_raddr     => ic_raddr,
         ic_rreq      => ic_rreq,
         io_dev       => io_dev,
         io_ix        => io_ix,
         io_mode      => io_mode,
         io_wdata     => io_wdata
      );
   uart_if_i : uart
      GENERIC MAP (
         baud            => 1_000_000,
         clock_frequency => 50_000_000
      )
      PORT MAP (
         clock               => clk,
         res_n               => res_n,
         data_stream_in      => data_stream_in,
         data_stream_in_stb  => data_stream_in_stb,
         data_stream_in_ack  => data_stream_in_ack,
         data_stream_in_done => data_stream_in_done,
         data_stream_out     => data_stream_out,
         data_stream_out_stb => data_stream_out_stb,
         tx                  => tx,
         rx                  => rx
      );

END struct;
