-- VHDL Entity riscvio_lib.obj_init_fsm.interface
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY riscvio_lib;
USE riscvio_lib.isa.all;
LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY obj_init_fsm IS
   PORT( 
      clk            : IN     std_logic;
      end_addr       : IN     word_T;
      pgu_mode_ex    : IN     pgu_mode_T;
      res_ex         : IN     reg_mem_T;
      res_n          : IN     std_logic;
      obj_init_addr  : OUT    word_T;
      obj_init_data  : OUT    word_T;
      obj_init_stall : OUT    boolean;
      obj_init_wr    : OUT    boolean
   );

-- Declarations

END obj_init_fsm ;
