-- VHDL Entity riscvio_lib.at_reg.interface
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY riscvio_lib;
USE riscvio_lib.isa.all;
LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY at_reg IS
   PORT( 
      clk            : IN     std_logic;
      ctrl_me        : IN     ctrl_sig_T;
      imm_me         : IN     word_T;
      obj_init_stall : IN     boolean;
      raux_me        : IN     raux_T;
      rdat_me        : IN     rdat_T;
      rdst_ix_me     : IN     reg_ix_T;
      res_at_u       : IN     reg_mem_T;
      res_n          : IN     std_logic;
      rptr_me        : IN     rptr_T;
      allocating_wb  : OUT    boolean;
      rd_wb          : OUT    reg_wb_T;
      rdst_ix_at     : OUT    reg_ix_T;
      res_at         : OUT    reg_mem_T
   );

-- Declarations

END at_reg ;
