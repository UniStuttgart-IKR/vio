-- VHDL Entity riscvio_lib.ex_reg.interface
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY riscvio_lib;
USE riscvio_lib.isa.all;
LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY ex_reg IS
   PORT( 
      clk                           : IN     std_logic;
      ctrl_dc                       : IN     ctrl_sig_T;
      frame_type_exception          : IN     boolean;
      imm_dc                        : IN     word_T;
      index_out_of_bounds_exception : IN     boolean;
      obj_init_stall                : IN     boolean;
      raux_dc                       : IN     raux_T;
      rdat_dc                       : IN     rdat_T;
      rdst_ix_dc                    : IN     reg_ix_T;
      res_ex_u                      : IN     reg_mem_T;
      res_n                         : IN     std_logic;
      rptr_dc                       : IN     rptr_T;
      state_error_dbu               : IN     boolean;
      state_error_pgu               : IN     boolean;
      allocating_me                 : OUT    boolean;
      ctrl_ex                       : OUT    ctrl_sig_T;
      imm_ex_reg                    : OUT    word_T;
      me_mode_dc_uq                 : OUT    mem_mode_t;
      me_mode_ex                    : OUT    mem_mode_T;
      pgu_mode_ex                   : OUT    pgu_mode_T;
      raux_dc_uq                    : OUT    raux_T;
      raux_ex_reg                   : OUT    raux_T;
      rdat_ex_reg                   : OUT    rdat_T;
      rdst_ix_ex_reg                : OUT    reg_ix_T;
      res_ex                        : OUT    reg_mem_T;
      res_ex_uq                     : OUT    reg_mem_T;
      rptr_dc_uq                    : OUT    rptr_T;
      rptr_ex_reg                   : OUT    rptr_T
   );

-- Declarations

END ex_reg ;
