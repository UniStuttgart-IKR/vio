--
-- VHDL Architecture riscvio_lib.alc_fwd_unit.behav
--
-- Created:
--          by - rbnlux.ckoehler (pc037)
--          at - 19:00:15 06/19/24
--
-- using Mentor Graphics HDL Designer(TM) 2022.3 Built on 14 Jul 2022 at 13:56:12
--
ARCHITECTURE behav OF alc_fwd_unit IS
BEGIN
END ARCHITECTURE behav;

