LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY riscvio_lib;
USE riscvio_lib.isa.all;
USE riscvio_lib.caches.all;
LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;
USE riscvio_lib.caches.all;

ENTITY me_res_mux IS
   PORT( 
      ctrl_ex      : IN     ctrl_sig_T;
      mem_out_me_u : IN     dword_T;
      raux_ex      : IN     raux_T;
      res_ex       : IN     reg_mem_T;
      res_me_u     : OUT    reg_mem_T
   );

-- Declarations

END me_res_mux ;
