--
-- VHDL Architecture riscvio_lib.block_ram_if.behav
--
-- Created:
--          by - rbnlux.ckoehler (pc038)
--          at - 16:10:55 06/05/24
--
-- using Mentor Graphics HDL Designer(TM) 2022.3 Built on 14 Jul 2022 at 13:56:12
--
ARCHITECTURE behav OF block_ram_if IS

BEGIN
--
--    -- read from RX Buffer 
--  read_p: process (all) is
--  begin  
--    -- assign default values
--    mem_out        <= (others => '0');
--    
--    if raddr_in_bounds then
--      case io_mode is
--        when lb =>
--          
--          case addr(1 downto 0) is
--            when "00" =>
--                rdata              <= (others => dcbr_data_a(BYTE0_RANGE'high));
--                mem_out(BYTE0_RANGE) <= dcbr_data_a(BYTE0_RANGE);
--                        
--            when "01" =>
--                rdata              <= (others => dcbr_data_a(BYTE1_RANGE'high));
--                mem_out(BYTE0_RANGE) <= dcbr_data_a(BYTE1_RANGE);
--                            
--            when "10" =>
--                rdata              <= (others => dcbr_data_a(BYTE2_RANGE'high));
--                mem_out(BYTE0_RANGE) <= dcbr_data_a(BYTE2_RANGE);
--                        
--            when "11" =>
--                rdata              <= (others => dcbr_data_a(BYTE3_RANGE'high));
--                mem_out(BYTE0_RANGE) <= dcbr_data_a(BYTE3_RANGE);
--            
--            when others =>
--                null;
--                
--          end case;
--          
--        when lbu =>
--          case addr(1 downto 0) is
--            when "00" =>
--                mem_out(BYTE0_RANGE) <= dcbr_data_a(BYTE0_RANGE); 
--                    
--            when "01" =>
--                mem_out(BYTE0_RANGE) <= dcbr_data_a(BYTE1_RANGE);
--                            
--            when "10" =>
--                mem_out(BYTE0_RANGE) <= dcbr_data_a(BYTE2_RANGE);
--                        
--            when "11" =>
--                mem_out(BYTE0_RANGE) <= dcbr_data_a(BYTE3_RANGE);
--                        
--            when others =>
--                null;
--                
--          end case;
--          
--        when lh =>
--          case addr(1) isdcbr_data_a
--            when "0" =>
--                rdata               <= (others => dcbr_data_a(HWORD0_RANGE'high));
--                mem_out(HWORD0_RANGE) <= dcbr_data_a(HWORD0_RANGE);
--                            
--            when "1" =>
--                rdata               <= (others => dcbr_data_a(HWORD1_RANGE'high));
--                mem_out(HWORD0_RANGE) <= dcbr_data_a(HWORD1_RANGE);
--                                
--            when others => 
--                null;
--            
--          end case;
--          
--        when lhu =>
--          case addr(1) is
--            when "0" =>
--                mem_out(HWORD0_RANGE) <= dcbr_data_a(HWORD0_RANGE);
--                            
--            when "1" =>
--                mem_out(HWORD0_RANGE) <= dcbr_data_a(HWORD1_RANGE);
--                            
--            when others => 
--                null;
--                
--          end case;
--  
--        when lw =>
--            mem_out <= dcbr_data_a;
--          
--        when others =>
--          null;
--      end case;
--    end if;
--  end process read_p;
--
--
--
--    -- write to IO Buffer
--  write_p: process (all) is
--  begin
--    -- assign default values
--    dcbr_byteena_a      <= (others => '0');
--    dcbr_data_a <= (others => '0');
--    dcbr_wren_a  <= '0';
--    
--    if waddr_in_bounds then
--      case io_mode is
--        when sb =>
--            dcbr_wren_a  <= '1';
--            byteena(to_integer(unsigned(addr(1 downto 0)))) <= '1';
--            wdata(BYTE0_RANGE) <= rdat.val(BYTE0_RANGE);
--            wdata(BYTE1_RANGE) <= rdat.val(BYTE0_RANGE);
--            wdata(BYTE2_RANGE) <= rdat.val(BYTE0_RANGE);
--            wdata(BYTE3_RANGE) <= rdat.val(BYTE0_RANGE);
--
--            
--        when sh =>
--            dcbr_wren_a  <= '1';
--            dcbr_byteena_a(to_integer(unsigned(addr(1) & '0'))) <= '1';
--            dcbr_byteena_a(to_integer(unsigned(addr(1) & '1'))) <= '1';
--            dcbr_data_a <= rdat.val(HWORD0_RANGE) 
--                             & rdat.val(HWORD0_RANGE) 
--               
--        when sw =>
--            dcbr_wren_a  <= '1';
--            dcbr_byteena_a <= X"F0" when addr(2) = '1' else X"0F";
--            dcbr_data_a <= rdat.val(WORD0_RANGE) & rdat.val(WORD0_RANGE);
--            
--        when sd =>
--          dcbr_wren_a  <= '1';
--          dcbr_byteena_a <= (others => '1');
--          dcbr_data_a <= rdat.val;
--  
--        when others =>
--          null;
--      end case;
--    end if;
--    
--  end process write_p;   
--
dram_wren_a  <= '0';
dram_byteena_a <= (others => '0');
END ARCHITECTURE behav;

