LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
LIBRARY riscvio_lib;
USE riscvio_lib.caches.all;
USE riscvio_lib.ISA.all;


ARCHITECTURE struct OF riscvio_tb IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL clk      : std_logic;
   SIGNAL ic_rack  : boolean;
   SIGNAL ic_raddr : std_logic_vector(ADDR_WIDTH - 1 DOWNTO 0) := (others => '0');
   SIGNAL ic_rdata : std_logic_vector(BUS_WIDTH - 1 DOWNTO 0);
   SIGNAL ic_rreq  : boolean                                   := false;
   SIGNAL res_n    : std_logic;


   -- Component Declarations
   COMPONENT clk_res_gen_var
   GENERIC (
      ONTIME    : time := 10 ns;
      OFFTIME   : time := 10 ns;
      RESETTIME : time := 35 ns
   );
   PORT (
      clk   : OUT    std_logic;
      res_n : OUT    std_logic
   );
   END COMPONENT;
   COMPONENT int_ram
   PORT (
      ac_raddr : IN     std_logic_vector (ADDR_WIDTH - 1 DOWNTO 0) := (others => '0');
      ac_rreq  : IN     boolean                                    := false;
      clk      : IN     std_logic;
      dc_raddr : IN     std_logic_vector (ADDR_WIDTH - 1 DOWNTO 0) := (others => '0');
      dc_rreq  : IN     boolean                                    := false;
      dc_waddr : IN     std_logic_vector (ADDR_WIDTH - 1 DOWNTO 0) := (others => '0');
      dc_wdata : IN     std_logic_vector (BUS_WIDTH - 1 DOWNTO 0)  := (others => '0');
      dc_wreq  : IN     boolean                                    := false;
      ic_raddr : IN     std_logic_vector (ADDR_WIDTH - 1 DOWNTO 0) := (others => '0');
      ic_rreq  : IN     boolean                                    := false;
      res_n    : IN     std_logic;
      ac_rack  : OUT    boolean;
      ac_rdata : OUT    std_logic_vector (BUS_WIDTH - 1 DOWNTO 0);
      dc_rack  : OUT    boolean;
      dc_rdata : OUT    std_logic_vector (BUS_WIDTH - 1 DOWNTO 0);
      dc_wack  : OUT    boolean;
      ic_rack  : OUT    boolean;
      ic_rdata : OUT    std_logic_vector (BUS_WIDTH - 1 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT riscvio
   PORT (
      clk      : IN     std_logic ;
      ic_rack  : IN     boolean ;
      ic_rdata : IN     std_logic_vector (BUS_WIDTH - 1 DOWNTO 0);
      res_n    : IN     std_logic ;
      ic_raddr : OUT    std_logic_vector (ADDR_WIDTH - 1 DOWNTO 0);
      ic_rreq  : OUT    boolean 
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : clk_res_gen_var USE ENTITY riscvio_lib.clk_res_gen_var;
   FOR ALL : int_ram USE ENTITY riscvio_lib.int_ram;
   FOR ALL : riscvio USE ENTITY riscvio_lib.riscvio;
   -- pragma synthesis_on


BEGIN

   -- Instance port mappings.
   clk_i : clk_res_gen_var
      GENERIC MAP (
         ONTIME    => 10 ns,
         OFFTIME   => 10 ns,
         RESETTIME => 35 ns
      )
      PORT MAP (
         clk   => clk,
         res_n => res_n
      );
   int_ram_i : int_ram
      PORT MAP (
         clk      => clk,
         res_n    => res_n,
         dc_rreq  => OPEN,
         dc_rack  => OPEN,
         dc_raddr => OPEN,
         dc_rdata => OPEN,
         ac_rreq  => OPEN,
         ac_rack  => OPEN,
         ac_raddr => OPEN,
         ac_rdata => OPEN,
         ic_rreq  => ic_rreq,
         ic_rack  => ic_rack,
         ic_raddr => ic_raddr,
         ic_rdata => ic_rdata,
         dc_wreq  => OPEN,
         dc_wack  => OPEN,
         dc_waddr => OPEN,
         dc_wdata => OPEN
      );
   riscvio_i : riscvio
      PORT MAP (
         clk      => clk,
         ic_rack  => ic_rack,
         ic_rdata => ic_rdata,
         res_n    => res_n,
         ic_raddr => ic_raddr,
         ic_rreq  => ic_rreq
      );

END struct;
