-- VHDL Architecture riscvio_lib.if_reg.behav
--
-- Created:
--          by - surfer.UNKNOWN (SURFER-A0000001)
--          at - 11:50:54 05.05.2024
--
-- using Mentor Graphics HDL Designer(TM) 2021.1 Built on 14 Jan 2021 at 15:11:42
--
ARCHITECTURE behav OF dc_reg IS
BEGIN
  process(clk, res_n) is
  begin
    if res_n = '0' then
      rdst_ix_dc_reg <= 0;
      rdat_dc_reg <= RDAT_NULL;
      rptr_dc_reg <= RPTR_NULL;
      raux_dc_reg <= RAUX_NULL;
      imm_dc_reg  <= (others => '0');
      ctrl_dc <= CTRL_NULL;
      pc_dc <= PC_NULL;
      branch_mode_dc <= no_branch;
      exc_dc <= well_behaved;
      ebreak_stall <= false;
    else
      if clk'event and clk = '1' then
        if pipe_flush then
          rdst_ix_dc_reg <= 0;
          rdat_dc_reg <= RDAT_NULL;
          rptr_dc_reg <= RPTR_NULL;
          raux_dc_reg <= RAUX_NULL;
          imm_dc_reg  <= (others => '0');
          ctrl_dc <= CTRL_NULL;
          pc_dc <= PC_NULL;
          branch_mode_dc <= no_branch;
          exc_dc <= well_behaved;
          ebreak_stall <= false;
        elsif not stall then
          if dbt_valid then
            ctrl_dc <= CTRL_NULL;
            branch_mode_dc <= no_branch;
            rdst_ix_dc_reg <= 0;
            rdat_dc_reg <= RDAT_NULL;
            rptr_dc_reg <= RPTR_NULL;
            raux_dc_reg <= RAUX_NULL;
            imm_dc_reg  <= (others => '0');
            exc_dc <= well_behaved;
            ebreak_stall <= false;
          else
            ctrl_dc <= ctrl_dc_u;
            branch_mode_dc <= ctrl_dc_u.branch_mode;
            rdst_ix_dc_reg <= rdst_ix_dc_u;
            rdat_dc_reg <= rdat_dc_u;
            rptr_dc_reg <= rptr_dc_u;
            raux_dc_reg <= raux_dc_u;
            imm_dc_reg  <= imm_dc_u;
            exc_dc <= exc_dc_u;
            ebreak_stall <= ctrl_dc_u.mnemonic = ebreak;
            --synthesis off
            assert ctrl_dc_u.mnemonic /= ebreak report "EBREAK" severity failure;
            --synthesis on
          end if;
          pc_dc <= pc_if;
        elsif ebreak_release then
          ebreak_stall <= false;
        end if;
      end if;
    end if;
  end process;

  alu_mode_dc     <= ctrl_dc.alu_mode; 
  alu_a_in_sel_dc <= ctrl_dc.alu_a_sel;
  alu_b_in_sel_dc <= ctrl_dc.alu_b_sel;
  res_mux_sel     <= ctrl_dc.ex_res_mux_sel;
  pgu_mode_dc     <= ctrl_dc.pgu_mode;
  fwd_allowed_dc  <= ctrl_dc.fwd_allowed;

END ARCHITECTURE behav;