LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY riscvio_lib;
USE riscvio_lib.isa.all;
USE riscvio_lib.pipeline.all;


ARCHITECTURE struct OF riscvio IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL REG_MEM_NULL_SIG   : reg_mem_T;
   SIGNAL a                  : word_T;
   SIGNAL ac_stall           : boolean;
   SIGNAL addr_me            : reg_mem_T;
   SIGNAL addr_me_uq         : reg_mem_T;
   SIGNAL allocating_at      : boolean;
   SIGNAL allocating_me      : boolean   := false;
   SIGNAL allocating_wb      : boolean;
   SIGNAL alu_a_in_sel_dc    : alu_in_sel_T;
   SIGNAL alu_b_in_sel_dc    : alu_in_sel_T;
   SIGNAL alu_mode_dc        : alu_mode_T;
   SIGNAL alu_out_ex_u       : word_T;
   SIGNAL at_mode            : at_mode_T;
   SIGNAL atomic_swap        : boolean;
   SIGNAL b                  : word_T;
   SIGNAL branch_mode_dc     : branch_mode_T;
   SIGNAL cjt                : pc_T;
   SIGNAL cjt_valid          : boolean;
   SIGNAL csr_ix             : reg_nbr_T;
   SIGNAL csr_mux_sel        : csr_mux_sel_T;
   SIGNAL csr_nbr            : reg_nbr_T;
   SIGNAL csr_reg            : reg_mem_T;
   SIGNAL ctrl_dc            : ctrl_sig_T;
   SIGNAL ctrl_dc_dec        : ctrl_sig_t;
   SIGNAL ctrl_dc_u          : ctrl_sig_T;
   SIGNAL ctrl_ex            : ctrl_sig_T;
   SIGNAL ctrl_me            : ctrl_sig_T;
   SIGNAL current_pc_d       : pc_T;
   SIGNAL current_pc_uq      : pc_T;
   SIGNAL dbt                : pc_T;
   SIGNAL dbt_valid          : boolean;
   SIGNAL dbu_exc            : exc_cause_T;
   SIGNAL dbu_out_ex_u       : reg_mem_T;
   SIGNAL dc_stall           : boolean;
   SIGNAL dt_at_u            : word_T;
   SIGNAL end_addr           : word_T;
   SIGNAL exc_dc             : exc_cause_T;
   SIGNAL exc_dc_dec         : exc_cause_T;
   SIGNAL exc_dc_u           : exc_cause_T;
   SIGNAL exc_ex             : exc_cause_T;
   SIGNAL exc_ex_u           : exc_cause_T;
   SIGNAL exc_me             : exc_cause_T;
   SIGNAL exc_wb             : exc_cause_T;
   SIGNAL false_sig          : boolean;
   SIGNAL flags              : alu_flags_T;
   SIGNAL fwd_allowed_dc     : boolean;
   SIGNAL fwd_allowed_ex     : boolean;
   SIGNAL ic_stall           : boolean;
   SIGNAL if_instr           : word_T;
   SIGNAL if_instr_d         : word_T;
   SIGNAL imm_dc             : word_T;
   SIGNAL imm_dc_reg         : word_T;
   SIGNAL imm_dc_u           : word_T;
   SIGNAL imm_dec            : word_T;
   SIGNAL imm_ex             : word_T;
   SIGNAL imm_ex_reg         : word_T;
   SIGNAL imm_me             : word_T;
   SIGNAL incremented_pc     : pc_T;
   SIGNAL insert_atomic      : boolean;
   SIGNAL insert_nop         : boolean;
   SIGNAL io_out_me_u        : word_T;
   SIGNAL io_stall_int       : boolean;
   SIGNAL me_addr            : mem_addr_T;
   SIGNAL me_addr_u          : mem_addr_T;
   SIGNAL me_addr_uq         : mem_addr_T;
   SIGNAL me_mode_ex         : mem_mode_T;
   SIGNAL me_mode_ex_uq      : mem_mode_T;
   SIGNAL mem_out_me_u       : dword_T;
   SIGNAL mux_exc            : exc_cause_T;
   SIGNAL next_obj_init_addr : word_T;
   SIGNAL obj_init_addr      : word_T;
   SIGNAL obj_init_byte_ena  : std_logic_vector(BUS_WIDTH/8 - 1 DOWNTO 0);
   SIGNAL obj_init_data      : buzz_word_T;
   SIGNAL obj_init_stall     : boolean;
   SIGNAL obj_init_wr        : boolean;
   SIGNAL pc_current_pc      : pc_T;
   SIGNAL pc_dc              : pc_T;
   SIGNAL pc_ex              : pc_T;
   SIGNAL pc_if              : pc_T;
   SIGNAL pc_me              : pc_T;
   SIGNAL pc_wb              : pc_T;
   SIGNAL pgu_exc            : exc_cause_T;
   SIGNAL pgu_mode_dc        : pgu_mode_T;
   SIGNAL pgu_mode_dc_uq     : pgu_mode_T;
   SIGNAL pgu_mode_ex        : pgu_mode_T;
   SIGNAL pgu_ptr_ex_u       : reg_mem_T;
   SIGNAL pi_at_u            : word_T;
   SIGNAL pipe_flush         : boolean;
   SIGNAL raux_dc            : raux_T;
   SIGNAL raux_dc_reg        : raux_T;
   SIGNAL raux_dc_u          : raux_T;
   SIGNAL raux_ex            : raux_T;
   SIGNAL raux_ex_reg        : raux_T;
   SIGNAL raux_ix            : reg_nbr_T;
   SIGNAL raux_me            : raux_T;
   SIGNAL raux_rf            : raux_T;
   SIGNAL rd_wb              : reg_wb_T;
   SIGNAL rdat_dc            : rdat_T;
   SIGNAL rdat_dc_reg        : rdat_T;
   SIGNAL rdat_dc_u          : rdat_T;
   SIGNAL rdat_ex            : rdat_T;
   SIGNAL rdat_ex_reg        : rdat_T;
   SIGNAL rdat_ix            : reg_nbr_T;
   SIGNAL rdat_me            : rdat_T;
   SIGNAL rdat_rf            : rdat_T;
   SIGNAL rdst_ix_at         : reg_nbr_T;
   SIGNAL rdst_ix_dc         : reg_nbr_T;
   SIGNAL rdst_ix_dc_reg     : reg_nbr_T;
   SIGNAL rdst_ix_dc_u       : reg_nbr_T;
   SIGNAL rdst_ix_dec        : reg_nbr_T;
   SIGNAL rdst_ix_ex         : reg_nbr_T;
   SIGNAL rdst_ix_ex_reg     : reg_nbr_T;
   SIGNAL rdst_ix_me         : reg_nbr_T := 0;
   SIGNAL res_at             : reg_mem_T;
   SIGNAL res_at_u           : reg_mem_T;
   SIGNAL res_ex             : reg_mem_T;
   SIGNAL res_ex_u           : reg_mem_T;
   SIGNAL res_me             : reg_mem_T;
   SIGNAL res_me_u           : reg_mem_T;
   SIGNAL res_mux_sel        : ex_res_mux_sel_T;
   SIGNAL rptr_dc            : rptr_T;
   SIGNAL rptr_dc_reg        : rptr_T;
   SIGNAL rptr_dc_u          : rptr_T;
   SIGNAL rptr_ex            : rptr_T;
   SIGNAL rptr_ex_reg        : rptr_T;
   SIGNAL rptr_ix            : reg_nbr_T;
   SIGNAL rptr_me            : rptr_T;
   SIGNAL rptr_rf            : rptr_T;
   SIGNAL sbt                : pc_T;
   SIGNAL sbt_valid          : boolean;
   SIGNAL stall              : boolean;
   SIGNAL start_addr         : word_T;
   SIGNAL start_addr_uq      : word_T;
   SIGNAL wdt_me             : word_T;
   SIGNAL wpi_me             : word_T;
   SIGNAL xret               : xret_T;
   SIGNAL zero_reg_ix        : reg_nbr_T := 0;


   -- Component Declarations
   COMPONENT ac_wrapper
   PORT (
      addr      : IN     reg_mem_T ;
      at_mode   : IN     at_mode_T ;
      clk       : IN     std_logic ;
      next_addr : IN     reg_mem_T ;
      rack      : IN     boolean ;
      rdata     : IN     buzz_word_T ;
      res_n     : IN     std_logic ;
      wack      : IN     boolean ;
      wdt       : IN     word_T ;
      wpi       : IN     word_T ;
      ldt       : OUT    word_T ;
      lpi       : OUT    word_T ;
      raddr     : OUT    std_logic_vector (31 DOWNTO 0);
      rreq      : OUT    boolean ;
      stall     : OUT    boolean ;
      waddr     : OUT    word_T ;
      wbyte_ena : OUT    std_logic_vector (BUS_WIDTH/8 - 1 DOWNTO 0);
      wdata     : OUT    buzz_word_T ;
      wreq      : OUT    boolean 
   );
   END COMPONENT;
   COMPONENT alu
   PORT (
      a       : IN     word_T ;
      b       : IN     word_T ;
      mode    : IN     alu_mode_T ;
      alu_out : OUT    word_T ;
      flags   : OUT    alu_flags_T 
   );
   END COMPONENT;
   COMPONENT alu_a_mux
   PORT (
      alu_a_in_sel : IN     alu_in_sel_T ;
      raux_dc      : IN     raux_T ;
      rdat_dc      : IN     rdat_T ;
      rptr_dc      : IN     rptr_T ;
      a            : OUT    word_T 
   );
   END COMPONENT;
   COMPONENT alu_b_mux
   PORT (
      alu_b_in_sel : IN     alu_in_sel_T ;
      imm_dc       : IN     word_T ;
      raux_dc      : IN     raux_T ;
      rdat_dc      : IN     rdat_T ;
      rptr_dc      : IN     rptr_T ;
      b            : OUT    word_T 
   );
   END COMPONENT;
   COMPONENT at_reg
   PORT (
      clk           : IN     std_logic ;
      ctrl_me       : IN     ctrl_sig_T ;
      exc_me        : IN     exc_cause_T ;
      imm_me        : IN     word_T ;
      pc_me         : IN     pc_T ;
      raux_me       : IN     raux_T ;
      rdat_me       : IN     rdat_T ;
      rdst_ix_me    : IN     reg_nbr_T ;
      res_at_u      : IN     reg_mem_T ;
      res_n         : IN     std_logic ;
      rptr_me       : IN     rptr_T ;
      stall         : IN     boolean ;
      allocating_wb : OUT    boolean ;
      exc_wb        : OUT    exc_cause_T ;
      pc_wb         : OUT    pc_T ;
      pipe_flush    : OUT    boolean ;
      rd_wb         : OUT    reg_wb_T ;
      rdst_ix_at    : OUT    reg_nbr_T ;
      res_at        : OUT    reg_mem_T 
   );
   END COMPONENT;
   COMPONENT at_res_mux
   PORT (
      ctrl_me  : IN     ctrl_sig_T ;
      dt_at_u  : IN     word_T ;
      pi_at_u  : IN     word_T ;
      res_me   : IN     reg_mem_T ;
      res_at_u : OUT    reg_mem_T 
   );
   END COMPONENT;
   COMPONENT clr_ptr_end_addr_mux
   PORT (
      raux_ex    : IN     raux_T ;
      rdst_ix_ex : IN     reg_nbr_T ;
      rptr_ex    : IN     rptr_T ;
      end_addr   : OUT    word_T 
   );
   END COMPONENT;
   COMPONENT csr_rf_mux
   PORT (
      csr_mux_sel : IN     csr_mux_sel_T ;
      csr_nbr     : IN     reg_nbr_T ;
      csr_reg     : IN     reg_mem_T ;
      raux_rf     : IN     raux_T ;
      rdat_rf     : IN     rdat_T ;
      rptr_rf     : IN     rptr_T ;
      raux_dc_u   : OUT    raux_T ;
      rdat_dc_u   : OUT    rdat_T ;
      rptr_dc_u   : OUT    rptr_T 
   );
   END COMPONENT;
   COMPONENT csr_unit
   PORT (
      clk       : IN     std_logic ;
      csr_ix    : IN     reg_nbr_T ;
      exc_wb    : IN     exc_cause_T ;
      pc_wb     : IN     pc_T ;
      rd_wb     : IN     reg_wb_T ;
      res_n     : IN     std_logic ;
      xret      : IN     xret_T ;
      cjt       : OUT    pc_T ;
      cjt_valid : OUT    boolean ;
      csr_nbr   : OUT    reg_nbr_T ;
      csr_reg   : OUT    reg_mem_T 
   );
   END COMPONENT;
   COMPONENT dc_reg
   PORT (
      clk             : IN     std_logic ;
      ctrl_dc_u       : IN     ctrl_sig_T ;
      dbt_valid       : IN     boolean ;
      exc_dc_u        : IN     exc_cause_T ;
      imm_dc_u        : IN     word_T ;
      pc_if           : IN     pc_T ;
      pipe_flush      : IN     boolean ;
      raux_dc_u       : IN     raux_T ;
      rdat_dc_u       : IN     rdat_T ;
      rdst_ix_dc_u    : IN     reg_nbr_T ;
      res_n           : IN     std_logic ;
      rptr_dc_u       : IN     rptr_T ;
      stall           : IN     boolean ;
      alu_a_in_sel_dc : OUT    alu_in_sel_T ;
      alu_b_in_sel_dc : OUT    alu_in_sel_T ;
      alu_mode_dc     : OUT    alu_mode_T ;
      branch_mode_dc  : OUT    branch_mode_T ;
      ctrl_dc         : OUT    ctrl_sig_T ;
      exc_dc          : OUT    exc_cause_T ;
      fwd_allowed_dc  : OUT    boolean ;
      imm_dc_reg      : OUT    word_T ;
      pc_dc           : OUT    pc_T ;
      pgu_mode_dc     : OUT    pgu_mode_T ;
      raux_dc_reg     : OUT    raux_T ;
      rdat_dc_reg     : OUT    rdat_T ;
      rdst_ix_dc_reg  : OUT    reg_nbr_T ;
      res_mux_sel     : OUT    ex_res_mux_sel_T ;
      rptr_dc_reg     : OUT    rptr_T 
   );
   END COMPONENT;
   COMPONENT dc_wrapper
   PORT (
      addr               : IN     mem_addr_T ;
      clk                : IN     std_logic ;
      mode               : IN     mem_mode_T ;
      next_addr          : IN     mem_addr_T ;
      next_mode          : IN     mem_mode_T ;
      next_obj_init_addr : IN     word_T ;
      obj_init_addr      : IN     word_T ;
      obj_init_byte_ena  : IN     std_logic_vector (BUS_WIDTH/8 - 1 DOWNTO 0);
      obj_init_data      : IN     buzz_word_T ;
      obj_init_wr        : IN     boolean ;
      rack               : IN     boolean ;
      rdata              : IN     buzz_word_T ;
      res_n              : IN     std_logic ;
      sd_raux            : IN     raux_T ;
      sd_rdat            : IN     rdat_T ;
      sd_rptr            : IN     rptr_T ;
      wack               : IN     boolean ;
      ld                 : OUT    dword_T ;
      raddr              : OUT    std_logic_vector (31 DOWNTO 0);
      rreq               : OUT    boolean ;
      stall              : OUT    boolean ;
      waddr              : OUT    std_logic_vector (31 DOWNTO 0);
      wbyte_ena          : OUT    std_logic_vector (BUS_WIDTH/8 - 1 DOWNTO 0);
      wdata              : OUT    buzz_word_T ;
      wreq               : OUT    boolean 
   );
   END COMPONENT;
   COMPONENT decoder
   PORT (
      atomic_swap : IN     boolean;
      instruction : IN     word_T;
      pc          : IN     pc_T;
      csr_ix      : OUT    csr_nbr_T;
      csr_mux_sel : OUT    csr_mux_sel_T;
      ctr_sig     : OUT    ctrl_sig_t;
      exc         : OUT    exc_cause_T;
      imm         : OUT    word_T;
      raux_ix     : OUT    reg_nbr_T;
      rdat_ix     : OUT    reg_nbr_T;
      rdst_ix     : OUT    reg_nbr_T;
      rptr_ix     : OUT    reg_nbr_T;
      sbt         : OUT    pc_T;
      sbt_valid   : OUT    boolean;
      xret        : OUT    xret_T
   );
   END COMPONENT;
   COMPONENT dyn_branch_unit
   PORT (
      alu_flags   : IN     alu_flags_T;
      branch_mode : IN     branch_mode_T;
      imm         : IN     word_T;
      pc          : IN     pc_T;
      raux        : IN     raux_T;
      rdat        : IN     rdat_T;
      rdst_ix     : IN     reg_nbr_T;
      rptr        : IN     rptr_T;
      dbt         : OUT    pc_T;
      dbt_valid   : OUT    boolean;
      dbu_exc     : OUT    exc_cause_T;
      ra_out      : OUT    reg_mem_T
   );
   END COMPONENT;
   COMPONENT ex_exc_encoder
   PORT (
      dbu_exc  : IN     exc_cause_T;
      mux_exc  : IN     exc_cause_T;
      pgu_exc  : IN     exc_cause_T;
      prev_exc : IN     exc_cause_T;
      exc      : OUT    exc_cause_T
   );
   END COMPONENT;
   COMPONENT ex_reg
   PORT (
      clk            : IN     std_logic ;
      ctrl_dc        : IN     ctrl_sig_T ;
      exc_ex_u       : IN     exc_cause_T ;
      imm_dc         : IN     word_T ;
      me_addr_u      : IN     mem_addr_T ;
      pc_dc          : IN     pc_T ;
      pipe_flush     : IN     boolean ;
      raux_dc        : IN     raux_T ;
      rdat_dc        : IN     rdat_T ;
      rdst_ix_dc     : IN     reg_nbr_T ;
      res_ex_u       : IN     reg_mem_T ;
      res_n          : IN     std_logic ;
      rptr_dc        : IN     rptr_T ;
      stall          : IN     boolean ;
      allocating_me  : OUT    boolean ;
      ctrl_ex        : OUT    ctrl_sig_T ;
      exc_ex         : OUT    exc_cause_T ;
      fwd_allowed_ex : OUT    boolean ;
      imm_ex_reg     : OUT    word_T ;
      me_addr        : OUT    mem_addr_T ;
      me_addr_uq     : OUT    mem_addr_T ;
      me_mode_ex     : OUT    mem_mode_T ;
      me_mode_ex_uq  : OUT    mem_mode_T ;
      pc_ex          : OUT    pc_T ;
      pgu_mode_dc_uq : OUT    pgu_mode_T ;
      pgu_mode_ex    : OUT    pgu_mode_T ;
      raux_ex_reg    : OUT    raux_T ;
      rdat_ex_reg    : OUT    rdat_T ;
      rdst_ix_ex_reg : OUT    reg_nbr_T ;
      res_ex         : OUT    reg_mem_T ;
      rptr_ex_reg    : OUT    rptr_T ;
      start_addr     : OUT    word_T ;
      start_addr_uq  : OUT    word_T 
   );
   END COMPONENT;
   COMPONENT ex_res_mux
   PORT (
      alu_mode_dc  : IN     alu_mode_T ;
      alu_out_ex_u : IN     word_T ;
      dbu_out_ex_u : IN     reg_mem_T ;
      pgu_ptr_ex_u : IN     reg_mem_T ;
      raux_dc      : IN     raux_T ;
      rdat_dc      : IN     rdat_T ;
      res_mux_sel  : IN     ex_res_mux_sel_T ;
      rptr_dc      : IN     rptr_T ;
      mux_exc      : OUT    exc_cause_T ;
      res_ex_u     : OUT    reg_mem_T 
   );
   END COMPONENT;
   COMPONENT fwd_unit
   PORT (
      fwd_0       : IN     boolean ;
      fwd_1       : IN     boolean ;
      fwd_2       : IN     boolean ;
      fwd_allowed : IN     boolean ;
      fwd_idx_0   : IN     reg_nbr_T  := 0;
      fwd_idx_1   : IN     reg_nbr_T  := 0;
      fwd_idx_2   : IN     reg_nbr_T  := 0;
      fwd_res_0   : IN     reg_mem_T  := REG_MEM_NULL;
      fwd_res_1   : IN     reg_mem_T  := REG_MEM_NULL;
      fwd_res_2   : IN     reg_mem_T  := REG_MEM_NULL;
      imm_reg     : IN     word_T ;
      raux_reg    : IN     raux_T ;
      rdat_reg    : IN     rdat_T ;
      rdst_reg    : IN     reg_nbr_T ;
      rptr_reg    : IN     rptr_T ;
      imm_fwd     : OUT    word_T ;
      raux_fwd    : OUT    raux_T ;
      rdat_fwd    : OUT    rdat_T ;
      rdst_fwd    : OUT    reg_nbr_T ;
      rptr_fwd    : OUT    rptr_T 
   );
   END COMPONENT;
   COMPONENT ic_wrapper
   PORT (
      clk        : IN     STD_LOGIC  := '1';
      dbranch    : IN     boolean;
      ic_rack    : IN     boolean;
      ic_rdata   : IN     std_logic_vector (BUS_WIDTH - 1 DOWNTO 0);
      next_pc    : IN     pc_T;
      pc         : IN     pc_T;
      pipe_flush : IN     boolean;
      res_n      : IN     std_logic;
      sbranch    : IN     boolean;
      ic_raddr   : OUT    std_logic_vector (ADDR_WIDTH - 1 DOWNTO 0);
      ic_rreq    : OUT    boolean;
      instr      : OUT    STD_LOGIC_VECTOR (31 DOWNTO 0);
      stall      : OUT    boolean
   );
   END COMPONENT;
   COMPONENT if_reg
   PORT (
      cjt_valid     : IN     boolean ;
      clk           : IN     std_logic ;
      dbt_valid     : IN     boolean ;
      if_instr_d    : IN     word_T ;
      insert_nop    : IN     boolean ;
      pc_current_pc : IN     pc_T ;
      pipe_flush    : IN     boolean ;
      res_n         : IN     std_logic ;
      sbt_valid     : IN     boolean ;
      stall         : IN     boolean ;
      if_instr      : OUT    word_T ;
      pc_if         : OUT    pc_T 
   );
   END COMPONENT;
   COMPONENT io_interface
   PORT (
      addr      : IN     mem_addr_T;
      io_rdata  : IN     word_T;
      io_stall  : IN     std_logic;
      mode      : IN     mem_mode_T;
      next_addr : IN     mem_addr_T;
      next_mode : IN     mem_mode_T;
      sd_raux   : IN     raux_T;
      sd_rdat   : IN     rdat_T;
      sd_rptr   : IN     rptr_T;
      io_dev    : OUT    std_logic_vector (11 DOWNTO 0);
      io_ix     : OUT    word_T;
      io_mode   : OUT    mem_mode_T;
      io_wdata  : OUT    word_T;
      ld        : OUT    word_T;
      stall     : OUT    boolean
   );
   END COMPONENT;
   COMPONENT me_reg
   PORT (
      clk           : IN     std_logic ;
      ctrl_ex       : IN     ctrl_sig_T ;
      exc_ex        : IN     exc_cause_T ;
      imm_ex        : IN     word_T ;
      pc_ex         : IN     pc_T ;
      pipe_flush    : IN     boolean ;
      raux_ex       : IN     raux_T ;
      rdat_ex       : IN     rdat_T ;
      rdst_ix_ex    : IN     reg_nbr_T ;
      res_me_u      : IN     reg_mem_T ;
      res_n         : IN     std_logic ;
      rptr_ex       : IN     rptr_T ;
      stall         : IN     boolean ;
      addr_me       : OUT    reg_mem_T ;
      addr_me_uq    : OUT    reg_mem_T ;
      allocating_at : OUT    boolean ;
      at_mode       : OUT    at_mode_T ;
      ctrl_me       : OUT    ctrl_sig_T ;
      exc_me        : OUT    exc_cause_T ;
      imm_me        : OUT    word_T ;
      pc_me         : OUT    pc_T ;
      raux_me       : OUT    raux_T ;
      rdat_me       : OUT    rdat_T ;
      rdst_ix_me    : OUT    reg_nbr_T ;
      res_me        : OUT    reg_mem_T ;
      rptr_me       : OUT    rptr_T ;
      wdt_me        : OUT    word_T ;
      wpi_me        : OUT    word_T 
   );
   END COMPONENT;
   COMPONENT me_res_mux
   PORT (
      ctrl_ex      : IN     ctrl_sig_T ;
      io_out_me_u  : IN     word_T ;
      mem_out_me_u : IN     dword_T ;
      raux_ex      : IN     raux_T ;
      res_ex       : IN     reg_mem_T ;
      rptr_ex      : IN     rptr_T ;
      res_me_u     : OUT    reg_mem_T 
   );
   END COMPONENT;
   COMPONENT next_pc_mux
   PORT (
      csr_pc            : IN     pc_T;
      csr_pc_valid      : IN     boolean;
      dbta_valid        : IN     boolean;
      dynamic_branch_pc : IN     pc_T;
      incremented_pc    : IN     pc_T;
      sbta_valid        : IN     boolean;
      static_branch_pc  : IN     pc_T;
      next_pc           : OUT    pc_T
   );
   END COMPONENT;
   COMPONENT nop_gen
   PORT (
      ctrl_dc_dec   : IN     ctrl_sig_t;
      exc_dc_dec    : IN     exc_cause_T;
      imm_dec       : IN     word_T;
      insert_atomic : IN     boolean;
      insert_nop    : IN     boolean;
      rdst_ix_dec   : IN     reg_nbr_T;
      ctrl_dc_u     : OUT    ctrl_sig_T;
      exc_dc_u      : OUT    exc_cause_T;
      imm_dc_u      : OUT    word_T;
      rdst_ix_dc_u  : OUT    reg_nbr_T
   );
   END COMPONENT;
   COMPONENT obj_init_fsm
   PORT (
      clk                : IN     std_logic ;
      dc_stall           : IN     boolean ;
      end_addr           : IN     word_T ;
      pgu_mode_dc_uq     : IN     pgu_mode_T ;
      pgu_mode_ex        : IN     pgu_mode_T ;
      rdst_ix_ex         : IN     reg_nbr_T ;
      res_n              : IN     std_logic ;
      start_addr         : IN     word_T ;
      start_addr_uq      : IN     word_T ;
      obj_init_byte_ena  : OUT    std_logic_vector (BUS_WIDTH/8 - 1 DOWNTO 0);
      obj_init_data      : OUT    buzz_word_T ;
      obj_init_stall     : OUT    boolean ;
      obj_init_wr        : OUT    boolean ;
      next_obj_init_addr : INOUT  word_T ;
      obj_init_addr      : INOUT  word_T 
   );
   END COMPONENT;
   COMPONENT pc_incrementer
   PORT (
      pc      : IN     pc_T;
      next_pc : OUT    pc_T
   );
   END COMPONENT;
   COMPONENT pc_reg
   PORT (
      cjt_valid     : IN     boolean ;
      clk           : IN     std_logic ;
      current_pc_d  : IN     pc_T ;
      dbt_valid     : IN     boolean ;
      insert_nop    : IN     boolean ;
      pipe_flush    : IN     boolean ;
      res_n         : IN     std_logic ;
      sbt_valid     : IN     boolean ;
      stall         : IN     boolean ;
      current_pc_uq : OUT    pc_T ;
      pc_current_pc : OUT    pc_T 
   );
   END COMPONENT;
   COMPONENT pgu
   PORT (
      imm      : IN     word_T ;
      pc       : IN     pc_T ;
      pgu_mode : IN     pgu_mode_T ;
      raux     : IN     raux_T ;
      rdat     : IN     rdat_T ;
      rdst_ix  : IN     reg_nbr_T ;
      rptr     : IN     rptr_T ;
      me_addr  : OUT    mem_addr_T ;
      pgu_exc  : OUT    exc_cause_T ;
      ptr      : OUT    reg_mem_T 
   );
   END COMPONENT;
   COMPONENT ral_nop_unit
   PORT (
      ctrl_dc       : IN     ctrl_sig_T;
      ctrl_ex       : IN     ctrl_sig_T;
      ctrl_if       : IN     ctrl_sig_T;
      dbt_valid     : IN     boolean;
      raux_ix       : IN     reg_nbr_T;
      rdat_ix       : IN     reg_nbr_T;
      rdst_dc       : IN     reg_nbr_T;
      rdst_ex       : IN     reg_nbr_T;
      rptr_ix       : IN     reg_nbr_T;
      sbt_valid     : IN     boolean;
      atomic_swap   : OUT    boolean;
      insert_atomic : OUT    boolean;
      insert_nop    : OUT    boolean
   );
   END COMPONENT;
   COMPONENT register_file
   PORT (
      clk     : IN     std_logic;
      raux_ix : IN     reg_nbr_T;
      rd_wb   : IN     reg_wb_T;
      rdat_ix : IN     reg_nbr_T;
      res_n   : IN     std_logic;
      rptr_ix : IN     reg_nbr_T;
      raux    : OUT    raux_T;
      rdat    : OUT    rdat_T;
      rptr    : OUT    rptr_T
   );
   END COMPONENT;
   COMPONENT stall_logic
   PORT (
      ac_stall       : IN     boolean ;
      clk            : IN     std_logic ;
      dc_stall       : IN     boolean ;
      ic_stall       : IN     boolean ;
      io_stall_int   : IN     boolean ;
      obj_init_stall : IN     boolean ;
      res_n          : IN     std_logic ;
      stall          : OUT    boolean 
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : ac_wrapper USE ENTITY riscvio_lib.ac_wrapper;
   FOR ALL : alu USE ENTITY riscvio_lib.alu;
   FOR ALL : alu_a_mux USE ENTITY riscvio_lib.alu_a_mux;
   FOR ALL : alu_b_mux USE ENTITY riscvio_lib.alu_b_mux;
   FOR ALL : at_reg USE ENTITY riscvio_lib.at_reg;
   FOR ALL : at_res_mux USE ENTITY riscvio_lib.at_res_mux;
   FOR ALL : clr_ptr_end_addr_mux USE ENTITY riscvio_lib.clr_ptr_end_addr_mux;
   FOR ALL : csr_rf_mux USE ENTITY riscvio_lib.csr_rf_mux;
   FOR ALL : csr_unit USE ENTITY riscvio_lib.csr_unit;
   FOR ALL : dc_reg USE ENTITY riscvio_lib.dc_reg;
   FOR ALL : dc_wrapper USE ENTITY riscvio_lib.dc_wrapper;
   FOR ALL : decoder USE ENTITY riscvio_lib.decoder;
   FOR ALL : dyn_branch_unit USE ENTITY riscvio_lib.dyn_branch_unit;
   FOR ALL : ex_exc_encoder USE ENTITY riscvio_lib.ex_exc_encoder;
   FOR ALL : ex_reg USE ENTITY riscvio_lib.ex_reg;
   FOR ALL : ex_res_mux USE ENTITY riscvio_lib.ex_res_mux;
   FOR ALL : fwd_unit USE ENTITY riscvio_lib.fwd_unit;
   FOR ALL : ic_wrapper USE ENTITY riscvio_lib.ic_wrapper;
   FOR ALL : if_reg USE ENTITY riscvio_lib.if_reg;
   FOR ALL : io_interface USE ENTITY riscvio_lib.io_interface;
   FOR ALL : me_reg USE ENTITY riscvio_lib.me_reg;
   FOR ALL : me_res_mux USE ENTITY riscvio_lib.me_res_mux;
   FOR ALL : next_pc_mux USE ENTITY riscvio_lib.next_pc_mux;
   FOR ALL : nop_gen USE ENTITY riscvio_lib.nop_gen;
   FOR ALL : obj_init_fsm USE ENTITY riscvio_lib.obj_init_fsm;
   FOR ALL : pc_incrementer USE ENTITY riscvio_lib.pc_incrementer;
   FOR ALL : pc_reg USE ENTITY riscvio_lib.pc_reg;
   FOR ALL : pgu USE ENTITY riscvio_lib.pgu;
   FOR ALL : ral_nop_unit USE ENTITY riscvio_lib.ral_nop_unit;
   FOR ALL : register_file USE ENTITY riscvio_lib.register_file;
   FOR ALL : stall_logic USE ENTITY riscvio_lib.stall_logic;
   -- pragma synthesis_on


BEGIN
   -- Architecture concurrent statements
   -- HDL Embedded Text Block 2 eb2
   -- eb2 2  
   REG_MEM_NULL_SIG <= REG_MEM_NULL;
   ZERO_REG_IX <= ali_T'pos(zero);       
   false_sig <= false;                              


   -- Instance port mappings.
   ac_i : ac_wrapper
      PORT MAP (
         addr      => addr_me,
         at_mode   => at_mode,
         clk       => clk,
         next_addr => addr_me_uq,
         rack      => ac_rack,
         rdata     => ac_rdata,
         res_n     => res_n,
         wack      => ac_wack,
         wdt       => wdt_me,
         wpi       => wpi_me,
         ldt       => pi_at_u,
         lpi       => dt_at_u,
         raddr     => ac_raddr,
         rreq      => ac_rreq,
         stall     => ac_stall,
         waddr     => ac_waddr,
         wbyte_ena => ac_wbyte_ena,
         wdata     => ac_wdata,
         wreq      => ac_wreq
      );
   alu_i : alu
      PORT MAP (
         a       => a,
         b       => b,
         mode    => alu_mode_dc,
         alu_out => alu_out_ex_u,
         flags   => flags
      );
   alu_a_mux_i : alu_a_mux
      PORT MAP (
         alu_a_in_sel => alu_a_in_sel_dc,
         raux_dc      => raux_dc,
         rdat_dc      => rdat_dc,
         rptr_dc      => rptr_dc,
         a            => a
      );
   alu_b_mux_i : alu_b_mux
      PORT MAP (
         alu_b_in_sel => alu_b_in_sel_dc,
         imm_dc       => imm_dc,
         raux_dc      => raux_dc,
         rdat_dc      => rdat_dc,
         rptr_dc      => rptr_dc,
         b            => b
      );
   at_reg_i : at_reg
      PORT MAP (
         clk           => clk,
         ctrl_me       => ctrl_me,
         exc_me        => exc_me,
         imm_me        => imm_me,
         pc_me         => pc_me,
         raux_me       => raux_me,
         rdat_me       => rdat_me,
         rdst_ix_me    => rdst_ix_me,
         res_at_u      => res_at_u,
         res_n         => res_n,
         rptr_me       => rptr_me,
         stall         => stall,
         allocating_wb => allocating_wb,
         exc_wb        => exc_wb,
         pc_wb         => pc_wb,
         pipe_flush    => pipe_flush,
         rd_wb         => rd_wb,
         rdst_ix_at    => rdst_ix_at,
         res_at        => res_at
      );
   at_res_mux_i : at_res_mux
      PORT MAP (
         ctrl_me  => ctrl_me,
         dt_at_u  => dt_at_u,
         pi_at_u  => pi_at_u,
         res_me   => res_me,
         res_at_u => res_at_u
      );
   clr_ptr_end_addr_mux_i : clr_ptr_end_addr_mux
      PORT MAP (
         raux_ex    => raux_ex,
         rdst_ix_ex => rdst_ix_ex,
         rptr_ex    => rptr_ex,
         end_addr   => end_addr
      );
   csr_rf_mux_i : csr_rf_mux
      PORT MAP (
         csr_mux_sel => csr_mux_sel,
         csr_nbr     => csr_nbr,
         csr_reg     => csr_reg,
         raux_rf     => raux_rf,
         rdat_rf     => rdat_rf,
         rptr_rf     => rptr_rf,
         raux_dc_u   => raux_dc_u,
         rdat_dc_u   => rdat_dc_u,
         rptr_dc_u   => rptr_dc_u
      );
   csr_unit_i : csr_unit
      PORT MAP (
         clk       => clk,
         csr_ix    => csr_ix,
         exc_wb    => exc_wb,
         pc_wb     => pc_wb,
         rd_wb     => rd_wb,
         res_n     => res_n,
         xret      => xret,
         cjt       => cjt,
         cjt_valid => cjt_valid,
         csr_nbr   => csr_nbr,
         csr_reg   => csr_reg
      );
   dc_reg_i : dc_reg
      PORT MAP (
         clk             => clk,
         ctrl_dc_u       => ctrl_dc_u,
         dbt_valid       => dbt_valid,
         exc_dc_u        => exc_dc_u,
         imm_dc_u        => imm_dc_u,
         pc_if           => pc_if,
         pipe_flush      => pipe_flush,
         raux_dc_u       => raux_dc_u,
         rdat_dc_u       => rdat_dc_u,
         rdst_ix_dc_u    => rdst_ix_dc_u,
         res_n           => res_n,
         rptr_dc_u       => rptr_dc_u,
         stall           => stall,
         alu_a_in_sel_dc => alu_a_in_sel_dc,
         alu_b_in_sel_dc => alu_b_in_sel_dc,
         alu_mode_dc     => alu_mode_dc,
         branch_mode_dc  => branch_mode_dc,
         ctrl_dc         => ctrl_dc,
         exc_dc          => exc_dc,
         fwd_allowed_dc  => fwd_allowed_dc,
         imm_dc_reg      => imm_dc_reg,
         pc_dc           => pc_dc,
         pgu_mode_dc     => pgu_mode_dc,
         raux_dc_reg     => raux_dc_reg,
         rdat_dc_reg     => rdat_dc_reg,
         rdst_ix_dc_reg  => rdst_ix_dc_reg,
         res_mux_sel     => res_mux_sel,
         rptr_dc_reg     => rptr_dc_reg
      );
   dc_i : dc_wrapper
      PORT MAP (
         addr               => me_addr,
         clk                => clk,
         mode               => me_mode_ex,
         next_addr          => me_addr_uq,
         next_mode          => me_mode_ex_uq,
         next_obj_init_addr => next_obj_init_addr,
         obj_init_addr      => obj_init_addr,
         obj_init_byte_ena  => obj_init_byte_ena,
         obj_init_data      => obj_init_data,
         obj_init_wr        => obj_init_wr,
         rack               => dc_rack,
         rdata              => dc_rdata,
         res_n              => res_n,
         sd_raux            => raux_ex,
         sd_rdat            => rdat_ex,
         sd_rptr            => rptr_ex,
         wack               => dc_wack,
         ld                 => mem_out_me_u,
         raddr              => dc_raddr,
         rreq               => dc_rreq,
         stall              => dc_stall,
         waddr              => dc_waddr,
         wbyte_ena          => dc_wbyte_ena,
         wdata              => dc_wdata,
         wreq               => dc_wreq
      );
   decoder_i : decoder
      PORT MAP (
         pc          => pc_if,
         instruction => if_instr,
         atomic_swap => atomic_swap,
         rdat_ix     => rdat_ix,
         rptr_ix     => rptr_ix,
         raux_ix     => raux_ix,
         csr_ix      => csr_ix,
         csr_mux_sel => csr_mux_sel,
         rdst_ix     => rdst_ix_dec,
         imm         => imm_dec,
         ctr_sig     => ctrl_dc_dec,
         sbt_valid   => sbt_valid,
         sbt         => sbt,
         exc         => exc_dc_dec,
         xret        => xret
      );
   dbu_i : dyn_branch_unit
      PORT MAP (
         rdat        => rdat_dc,
         raux        => raux_dc,
         rptr        => rptr_dc,
         imm         => imm_dc,
         rdst_ix     => rdst_ix_dc,
         alu_flags   => flags,
         branch_mode => branch_mode_dc,
         pc          => pc_dc,
         dbu_exc     => dbu_exc,
         ra_out      => dbu_out_ex_u,
         dbt_valid   => dbt_valid,
         dbt         => dbt
      );
   ex_exc_i : ex_exc_encoder
      PORT MAP (
         prev_exc => exc_dc,
         exc      => exc_ex_u,
         mux_exc  => mux_exc,
         dbu_exc  => dbu_exc,
         pgu_exc  => pgu_exc
      );
   ex_reg_i : ex_reg
      PORT MAP (
         clk            => clk,
         ctrl_dc        => ctrl_dc,
         exc_ex_u       => exc_ex_u,
         imm_dc         => imm_dc,
         me_addr_u      => me_addr_u,
         pc_dc          => pc_dc,
         pipe_flush     => pipe_flush,
         raux_dc        => raux_dc,
         rdat_dc        => rdat_dc,
         rdst_ix_dc     => rdst_ix_dc,
         res_ex_u       => res_ex_u,
         res_n          => res_n,
         rptr_dc        => rptr_dc,
         stall          => stall,
         allocating_me  => allocating_me,
         ctrl_ex        => ctrl_ex,
         exc_ex         => exc_ex,
         fwd_allowed_ex => fwd_allowed_ex,
         imm_ex_reg     => imm_ex_reg,
         me_addr        => me_addr,
         me_addr_uq     => me_addr_uq,
         me_mode_ex     => me_mode_ex,
         me_mode_ex_uq  => me_mode_ex_uq,
         pc_ex          => pc_ex,
         pgu_mode_dc_uq => pgu_mode_dc_uq,
         pgu_mode_ex    => pgu_mode_ex,
         raux_ex_reg    => raux_ex_reg,
         rdat_ex_reg    => rdat_ex_reg,
         rdst_ix_ex_reg => rdst_ix_ex_reg,
         res_ex         => res_ex,
         rptr_ex_reg    => rptr_ex_reg,
         start_addr     => start_addr,
         start_addr_uq  => start_addr_uq
      );
   ex_res_mux_i : ex_res_mux
      PORT MAP (
         alu_mode_dc  => alu_mode_dc,
         alu_out_ex_u => alu_out_ex_u,
         dbu_out_ex_u => dbu_out_ex_u,
         pgu_ptr_ex_u => pgu_ptr_ex_u,
         raux_dc      => raux_dc,
         rdat_dc      => rdat_dc,
         res_mux_sel  => res_mux_sel,
         rptr_dc      => rptr_dc,
         mux_exc      => mux_exc,
         res_ex_u     => res_ex_u
      );
   fwd_ex_i : fwd_unit
      PORT MAP (
         fwd_0       => allocating_me,
         fwd_1       => allocating_at,
         fwd_2       => allocating_wb,
         fwd_allowed => fwd_allowed_dc,
         fwd_idx_0   => rdst_ix_ex_reg,
         fwd_idx_1   => rdst_ix_me,
         fwd_idx_2   => rdst_ix_at,
         fwd_res_0   => res_ex,
         fwd_res_1   => res_me,
         fwd_res_2   => res_at,
         imm_reg     => imm_dc_reg,
         raux_reg    => raux_dc_reg,
         rdat_reg    => rdat_dc_reg,
         rdst_reg    => rdst_ix_dc_reg,
         rptr_reg    => rptr_dc_reg,
         imm_fwd     => imm_dc,
         raux_fwd    => raux_dc,
         rdat_fwd    => rdat_dc,
         rdst_fwd    => rdst_ix_dc,
         rptr_fwd    => rptr_dc
      );
   fwd_me_i : fwd_unit
      PORT MAP (
         fwd_0       => false_sig,
         fwd_1       => false_sig,
         fwd_2       => false_sig,
         fwd_allowed => fwd_allowed_ex,
         fwd_idx_0   => rdst_ix_me,
         fwd_idx_1   => zero_reg_ix,
         fwd_idx_2   => zero_reg_ix,
         fwd_res_0   => res_me,
         fwd_res_1   => res_at,
         fwd_res_2   => REG_MEM_NULL_SIG,
         imm_reg     => imm_ex_reg,
         raux_reg    => raux_ex_reg,
         rdat_reg    => rdat_ex_reg,
         rdst_reg    => rdst_ix_ex_reg,
         rptr_reg    => rptr_ex_reg,
         imm_fwd     => imm_ex,
         raux_fwd    => raux_ex,
         rdat_fwd    => rdat_ex,
         rdst_fwd    => rdst_ix_ex,
         rptr_fwd    => rptr_ex
      );
   ic_i : ic_wrapper
      PORT MAP (
         pc         => pc_current_pc,
         next_pc    => current_pc_uq,
         clk        => clk,
         res_n      => res_n,
         instr      => if_instr_d,
         stall      => ic_stall,
         sbranch    => sbt_valid,
         dbranch    => dbt_valid,
         pipe_flush => pipe_flush,
         ic_rreq    => ic_rreq,
         ic_rack    => ic_rack,
         ic_raddr   => ic_raddr,
         ic_rdata   => ic_rdata
      );
   if_reg_i : if_reg
      PORT MAP (
         cjt_valid     => cjt_valid,
         clk           => clk,
         dbt_valid     => dbt_valid,
         if_instr_d    => if_instr_d,
         insert_nop    => insert_nop,
         pc_current_pc => pc_current_pc,
         pipe_flush    => pipe_flush,
         res_n         => res_n,
         sbt_valid     => sbt_valid,
         stall         => stall,
         if_instr      => if_instr,
         pc_if         => pc_if
      );
   io_if_i : io_interface
      PORT MAP (
         addr      => me_addr,
         next_addr => me_addr_uq,
         sd_rdat   => rdat_ex,
         sd_rptr   => rptr_ex,
         sd_raux   => raux_ex,
         mode      => me_mode_ex,
         next_mode => me_mode_ex_uq,
         ld        => io_out_me_u,
         stall     => io_stall_int,
         io_wdata  => io_wdata,
         io_rdata  => io_rdata,
         io_ix     => io_ix,
         io_dev    => io_dev,
         io_mode   => io_mode,
         io_stall  => io_stall
      );
   me_reg_i : me_reg
      PORT MAP (
         clk           => clk,
         ctrl_ex       => ctrl_ex,
         exc_ex        => exc_ex,
         imm_ex        => imm_ex,
         pc_ex         => pc_ex,
         pipe_flush    => pipe_flush,
         raux_ex       => raux_ex,
         rdat_ex       => rdat_ex,
         rdst_ix_ex    => rdst_ix_ex,
         res_me_u      => res_me_u,
         res_n         => res_n,
         rptr_ex       => rptr_ex,
         stall         => stall,
         addr_me       => addr_me,
         addr_me_uq    => addr_me_uq,
         allocating_at => allocating_at,
         at_mode       => at_mode,
         ctrl_me       => ctrl_me,
         exc_me        => exc_me,
         imm_me        => imm_me,
         pc_me         => pc_me,
         raux_me       => raux_me,
         rdat_me       => rdat_me,
         rdst_ix_me    => rdst_ix_me,
         res_me        => res_me,
         rptr_me       => rptr_me,
         wdt_me        => wdt_me,
         wpi_me        => wpi_me
      );
   me_res_mux_i : me_res_mux
      PORT MAP (
         ctrl_ex      => ctrl_ex,
         io_out_me_u  => io_out_me_u,
         mem_out_me_u => mem_out_me_u,
         raux_ex      => raux_ex,
         res_ex       => res_ex,
         rptr_ex      => rptr_ex,
         res_me_u     => res_me_u
      );
   next_pc_mux_i : next_pc_mux
      PORT MAP (
         incremented_pc    => incremented_pc,
         static_branch_pc  => sbt,
         dynamic_branch_pc => dbt,
         csr_pc            => cjt,
         dbta_valid        => dbt_valid,
         sbta_valid        => sbt_valid,
         csr_pc_valid      => cjt_valid,
         next_pc           => current_pc_d
      );
   nop_gen_i : nop_gen
      PORT MAP (
         ctrl_dc_dec   => ctrl_dc_dec,
         ctrl_dc_u     => ctrl_dc_u,
         imm_dc_u      => imm_dc_u,
         imm_dec       => imm_dec,
         exc_dc_dec    => exc_dc_dec,
         exc_dc_u      => exc_dc_u,
         insert_nop    => insert_nop,
         insert_atomic => insert_atomic,
         rdst_ix_dc_u  => rdst_ix_dc_u,
         rdst_ix_dec   => rdst_ix_dec
      );
   obj_init_fsm_i : obj_init_fsm
      PORT MAP (
         clk                => clk,
         dc_stall           => dc_stall,
         end_addr           => end_addr,
         pgu_mode_dc_uq     => pgu_mode_dc_uq,
         pgu_mode_ex        => pgu_mode_ex,
         rdst_ix_ex         => rdst_ix_ex,
         res_n              => res_n,
         start_addr         => start_addr,
         start_addr_uq      => start_addr_uq,
         obj_init_byte_ena  => obj_init_byte_ena,
         obj_init_data      => obj_init_data,
         obj_init_stall     => obj_init_stall,
         obj_init_wr        => obj_init_wr,
         next_obj_init_addr => next_obj_init_addr,
         obj_init_addr      => obj_init_addr
      );
   pc_increment_i : pc_incrementer
      PORT MAP (
         pc      => pc_current_pc,
         next_pc => incremented_pc
      );
   pc_reg_i : pc_reg
      PORT MAP (
         cjt_valid     => cjt_valid,
         clk           => clk,
         current_pc_d  => current_pc_d,
         dbt_valid     => dbt_valid,
         insert_nop    => insert_nop,
         pipe_flush    => pipe_flush,
         res_n         => res_n,
         sbt_valid     => sbt_valid,
         stall         => stall,
         current_pc_uq => current_pc_uq,
         pc_current_pc => pc_current_pc
      );
   pgu_i : pgu
      PORT MAP (
         imm      => imm_dc,
         pc       => pc_dc,
         pgu_mode => pgu_mode_dc,
         raux     => raux_dc,
         rdat     => rdat_dc,
         rdst_ix  => rdst_ix_dc,
         rptr     => rptr_dc,
         me_addr  => me_addr_u,
         pgu_exc  => pgu_exc,
         ptr      => pgu_ptr_ex_u
      );
   ral_nop_i : ral_nop_unit
      PORT MAP (
         ctrl_if       => ctrl_dc_dec,
         ctrl_dc       => ctrl_dc,
         ctrl_ex       => ctrl_ex,
         rdat_ix       => rdat_ix,
         raux_ix       => raux_ix,
         rptr_ix       => rptr_ix,
         rdst_dc       => rdst_ix_dc,
         rdst_ex       => rdst_ix_ex,
         sbt_valid     => sbt_valid,
         dbt_valid     => dbt_valid,
         atomic_swap   => atomic_swap,
         insert_atomic => insert_atomic,
         insert_nop    => insert_nop
      );
   register_file_i : register_file
      PORT MAP (
         clk     => clk,
         res_n   => res_n,
         rdat_ix => rdat_ix,
         rptr_ix => rptr_ix,
         raux_ix => raux_ix,
         rdat    => rdat_rf,
         rptr    => rptr_rf,
         raux    => raux_rf,
         rd_wb   => rd_wb
      );
   stall_logic_i : stall_logic
      PORT MAP (
         ac_stall       => ac_stall,
         clk            => clk,
         dc_stall       => dc_stall,
         ic_stall       => ic_stall,
         io_stall_int   => io_stall_int,
         obj_init_stall => obj_init_stall,
         res_n          => res_n,
         stall          => stall
      );

END struct;
