--
-- VHDL Architecture riscvio_lib.dual_port_ram.mixed
--
-- Created:
--          by - rbnlux.ckoehler (pc037)
--          at - 15:00:43 05/15/24
--
-- using Mentor Graphics HDL Designer(TM) 2022.3 Built on 14 Jul 2022 at 13:56:12
--

LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY dualportram IS
	PORT
	(
		address_a		: IN STD_LOGIC_VECTOR (ADDR_W - 1 DOWNTO 0);
		address_b		: IN STD_LOGIC_VECTOR (ADDR_W - 1 DOWNTO 0);
		clock		: IN STD_LOGIC  := '1';
		data_a		: IN STD_LOGIC_VECTOR (DATAW - 1 DOWNTO 0);
		data_b		: IN STD_LOGIC_VECTOR (DATAW - 1 DOWNTO 0);
		wren_a		: IN STD_LOGIC  := '0';
		wren_b		: IN STD_LOGIC  := '0';
		q_a		    : OUT STD_LOGIC_VECTOR (DATAW - 1 DOWNTO 0);
		q_b		    : OUT STD_LOGIC_VECTOR (DATAW - 1 DOWNTO 0)
	);
END dualportram;

ARCHITECTURE mixed OF dual_port_ram IS
    SIGNAL sub_wire0	: STD_LOGIC_VECTOR (DATAW - 1 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (DATAW - 1 DOWNTO 0);
BEGIN
    q_a    <= sub_wire0;
	q_b    <= sub_wire1;

	altsyncram_component : altsyncram
	GENERIC MAP (
		address_reg_b => "CLOCK0",
		clock_enable_input_a => "BYPASS",
		clock_enable_input_b => "BYPASS",
		clock_enable_output_a => "BYPASS",
		clock_enable_output_b => "BYPASS",
		indata_reg_b => "CLOCK0",
		init_file => INIT_FILE,
		intended_device_family => "Cyclone V",
		lpm_type => "altsyncram",
		numwords_a => SIZE_WORDS,
		numwords_b => SIZE_WORDS,
		operation_mode => "BIDIR_DUAL_PORT",
		outdata_aclr_a => "NONE",
		outdata_aclr_b => "NONE",
		outdata_reg_a => "UNREGISTERED",
		outdata_reg_b => "UNREGISTERED",
		power_up_uninitialized => "FALSE",
		read_during_write_mode_mixed_ports => "DONT_CARE",
		read_during_write_mode_port_a => "NEW_DATA_NO_NBE_READ",
		read_during_write_mode_port_b => "NEW_DATA_NO_NBE_READ",
		widthad_a => ADDR_W,
		widthad_b => ADDR_W,
		width_a => DATAW,
		width_b => DATAW,
		width_byteena_a => 1,
		width_byteena_b => 1,
		wrcontrol_wraddress_reg_b => "CLOCK0"
	)
	PORT MAP (
		address_a => address_a,
		address_b => address_b,
		clock0 => clock,
		data_a => data_a,
		data_b => data_b,
		wren_a => wren_a,
		wren_b => wren_b,
		q_a => sub_wire0,
		q_b => sub_wire1
	);
END ARCHITECTURE mixed;

